library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package pkg is
    type slv8_array_t is array (natural range <>) of std_logic_vector(31 downto 0);
    type mem_array_t is array (natural range <>) of std_logic_vector(7 downto 0);
end package;

package body pkg is
end package body;