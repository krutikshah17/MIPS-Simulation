library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;
library work;
use work.pkg.all;


entity Data_Memory is
port (   clk_DM                  : in std_logic;
         reset_DM                : in std_logic;   
         mem_access_addr_DM      : in std_logic_Vector(31 downto 0);
         mem_write_data_DM       : in std_logic_Vector(31 downto 0);
         mem_write_en_DM         : in std_logic;
         mem_read_DM             : in std_logic;
         mem_read_data_DM        : out std_logic_Vector(31 downto 0);
         key_vld_DM              : in std_logic;
         ukey_DM                 : in std_logic_Vector(31 downto 0);
--         array_m                 : out mem_array_t(0 to 1023);

         
         din_DM                  : in  std_logic_vector(63 downto 0);
         di_vld_DM               : in std_logic;
         mode_DM                    : in std_logic_vector(3 downto 0)
     );
end Data_Memory;


architecture Behavioral of Data_Memory is

signal i: integer;
signal ram_addr  : std_logic_vector(7 downto 0);

type data_mem is array (0 to 1023 ) of std_logic_vector (7 downto 0); 
--signal RAM: mem_array_t(0 to 1023);

signal RAM: data_mem; 

--:= data_mem'(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--A,B --0-7 

--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--S0=0,S1=0 --8-15 
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--s2,s3 --16-23
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--s4,s5 --24-31
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--s6,s7 --32-39
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--s8,s9 --40-47
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--s10,s11 --48-55
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--s12,s13 --56-63
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--s14,s15 --64-71
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--s16,s17 --72-79
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--s18,s19 --80-87
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--s20,s21 --88-95
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--s22,s23  --96-103
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--s24,s25 --104-111
                                  
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--L[3],L[2] --112-119
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--L[1],L[0] --120-127
                                  
--                                  x"B7", x"E1", x"51", x"63", x"9E", x"37", x"79", x"B9",--P,Q --128-135
                                  
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--136-143 --mode,di_vld
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --144-151--key_vld,ukey
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--152-159
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --160-167
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --168-175
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --176-183
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --184-191
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --192-199
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --200-207
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --208-215
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --216-223
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --224-231
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --232-239
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --240-247
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --248-255
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--136-263
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --144-271
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--152-279
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --160-287
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --168-295
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --176-303
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --184-311
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --192-319
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --200-327
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --208-335
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --216-343
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --224-351
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --232-359
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --240-367
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --248-375
--                                        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--136-143
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --144-151
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--152-159
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --160-167
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --168-175
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --176-183
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --184-191
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --192-199
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --200-207
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --208-215
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --216-223
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --224-231
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --232-239
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --240-247
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --248-255
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--136-263
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --144-271
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--152-279
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --160-287
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --168-295
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --176-303
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --184-311
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --192-319
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --200-327
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --208-335
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --216-343
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --224-351
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --232-359
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --240-367
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --248-375
--                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--136-143
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --144-151
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--152-159
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --160-167
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --168-175
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --176-183
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --184-191
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --192-199
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --200-207
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --208-215
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --216-223
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --224-231
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --232-239
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --240-247
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --248-255
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--136-263
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --144-271
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--152-279
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --160-287
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --168-295
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --176-303
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --184-311
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --192-319
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --200-327
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --208-335
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --216-343
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --224-351
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --232-359
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --240-367
--                                          x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --248-375
--                                            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--136-143
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --144-151
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--152-159
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --160-167
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --168-175
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --176-183
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --184-191
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --192-199
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --200-207
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --208-215
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --216-223
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --224-231
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --232-239
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --240-247
--                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --248-255
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--136-263
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --144-271
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--152-279
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --160-287
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --168-295
--                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00" --1017-1023
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --184-311
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --192-319
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --200-327
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --208-335
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --216-343
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --224-351
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --232-359
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --240-367
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --248-375
----                                      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--136-143
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --144-151
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--152-159
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --160-167
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --168-175
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --176-183
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --184-191
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --192-199
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --200-207
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --208-215
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --216-223
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --224-231
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --232-239
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --240-247
----                                    x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --248-255
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--136-263
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --144-271
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",--152-279
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --160-287
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --168-295
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --176-303
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --184-311
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --192-319
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --200-327
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --208-335
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --216-343
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --224-351
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --232-359
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --240-367
----                                  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00" --248-1335
                                  
                                                                    
                                                                       
--                                  );

begin

 ram_addr <= mem_access_addr_DM(7 downto 0);

 process(key_vld_DM,ukey_DM, clk_DM, ram_addr, mem_write_en_DM, mem_write_data_DM,reset_DM)
 begin
 
 if(reset_DM = '1') then
 
     RAM(7) <= din_DM(7 downto 0);
     RAM(6) <= din_DM(15 downto 8);
     RAM(5) <= din_DM(23 downto 16);
     RAM(4) <= din_DM(31 downto 24);
     RAM(3) <= din_DM(39 downto 32);
     RAM(2) <= din_DM(47 downto 40);
     RAM(1) <= din_DM(55 downto 48);
     RAM(0) <= din_DM(63 downto 56);
             
     RAM(151) <= ukey_DM(7 downto 0);
     RAM(150) <= ukey_DM(15 downto 8);
     RAM(149) <= ukey_DM(23 downto 16);
     RAM(148) <= ukey_DM(31 downto 24);
     
      --Mode
     RAM(136) <= x"00";
     RAM(137) <= x"00";
     RAM(138) <= x"00";
     RAM(139) <= "00000000";
     
     --Di_Valid
     RAM(140) <= x"00";
     RAM(141) <= x"00";
     RAM(142) <= x"00";
     RAM(143) <= "00000000";
     
     --Key Valid
     RAM(144) <= x"00";
     RAM(145) <= x"00";
     RAM(146) <= x"00";
     RAM(147) <= "00000000";
     
--      --Mode
--      if (mode_DM = x"1" or mode_DM = x"2" or mode_DM = x"4" or mode_DM = x"8") then
--          RAM(136) <= x"00";
--          RAM(137) <= x"00";
--          RAM(138) <= x"00";
--          RAM(139) <= "0000" & mode_DM;
--      end if;

--     if (di_vld_DM = '1') then

            
----          --Mode
----          RAM(136) <= x"00";
----          RAM(137) <= x"00";
----          RAM(138) <= x"00";
----          RAM(139) <= "0000" & mode_DM;
          
--          --Di_Valid
--          RAM(140) <= x"00";
--          RAM(141) <= x"00";
--          RAM(142) <= x"00";
--          RAM(143) <= "0000000" & di_vld_DM;
          
--        --Key Valid
--         RAM(144) <= x"00";
--         RAM(145) <= x"00";
--         RAM(146) <= x"00";
--         RAM(147) <= "00000000";
                 
--     end if;  
 
     if (key_vld_DM = '1') then
        
     
    
         FOR i IN 8 TO 111 LOOP
             RAM(i)<=(OTHERS=>'0');
         END LOOP;
         
         FOR i IN 116 TO 127 LOOP
             RAM(i)<=(OTHERS=>'0');
         END LOOP;
         
         RAM(128) <= x"B7";
         RAM(129) <= x"E1"; 
         RAM(130) <= x"51"; 
         RAM(131) <= x"63"; 
         RAM(132) <= x"9E"; 
         RAM(133) <= x"37"; 
         RAM(134) <= x"79"; 
         RAM(135) <= x"B9";  
         
--         --Mode
--         RAM(136) <= x"00";
--         RAM(137) <= x"00";
--         RAM(138) <= x"00";
--         RAM(139) <= "00000000";
         
--         --Di_Valid
--         RAM(140) <= x"00";
--         RAM(141) <= x"00";
--         RAM(142) <= x"00";
--         RAM(143) <= "00000000";
         
--         --Key Valid
--         RAM(144) <= x"00";
--         RAM(145) <= x"00";
--         RAM(146) <= x"00";
--         RAM(147) <= "00000000";
         
         FOR i IN 148 TO 1023 LOOP
             RAM(i)<=(OTHERS=>'0');
         END LOOP;
    end if; 
    
 elsif(rising_edge(clk_DM)) then
 
     RAM(7) <= din_DM(7 downto 0);
     RAM(6) <= din_DM(15 downto 8);
     RAM(5) <= din_DM(23 downto 16);
     RAM(4) <= din_DM(31 downto 24);
     RAM(3) <= din_DM(39 downto 32);
     RAM(2) <= din_DM(47 downto 40);
     RAM(1) <= din_DM(55 downto 48);
     RAM(0) <= din_DM(63 downto 56);
     
     RAM(151) <= ukey_DM(7 downto 0);
     RAM(150) <= ukey_DM(15 downto 8);
     RAM(149) <= ukey_DM(23 downto 16);
     RAM(148) <= ukey_DM(31 downto 24);
     
--     if (mode_DM = x"1" or mode_DM = x"2" or mode_DM = x"4" or mode_DM = x"8") then
--        RAM(136) <= x"00";
--        RAM(137) <= x"00";
--        RAM(138) <= x"00";
--        RAM(139) <= "0000" & mode_DM;
--     end if;
         
    if (mem_write_en_DM='1') then
             ram(to_integer(unsigned(ram_addr)))   <= mem_write_data_DM(31 downto 24);
             ram(to_integer(unsigned(ram_addr)+1)) <= mem_write_data_DM(23 downto 16);
             ram(to_integer(unsigned(ram_addr)+2)) <= mem_write_data_DM(15 downto 8);
             ram(to_integer(unsigned(ram_addr)+3)) <= mem_write_data_DM(7 downto 0);
             
--     elsif (di_vld_DM = '1') then
--         RAM(7) <= din_DM(7 downto 0);
--         RAM(6) <= din_DM(15 downto 8);
--         RAM(5) <= din_DM(23 downto 16);
--         RAM(4) <= din_DM(31 downto 24);
--         RAM(3) <= din_DM(39 downto 32);
--         RAM(2) <= din_DM(47 downto 40);
--         RAM(1) <= din_DM(55 downto 48);
--         RAM(0) <= din_DM(63 downto 56);
         
         --Mode
--         RAM(136) <= x"00";
--         RAM(137) <= x"00";
--         RAM(138) <= x"00";
--         RAM(139) <= "0000" & mode_DM;
         
--         --Di_Valid
--         RAM(140) <= x"00";
--         RAM(141) <= x"00";
--         RAM(142) <= x"00";
--         RAM(143) <= "0000000" & di_vld_DM;
         
--       --Key Valid
--        RAM(144) <= x"00";
--        RAM(145) <= x"00";
--        RAM(146) <= x"00";
--        RAM(147) <= "00000000";
      
--      elsif (key_vld_DM = '1') then
--         RAM(115) <= ukey_DM(7 downto 0);
--         RAM(114) <= ukey_DM(15 downto 8);
--         RAM(113) <= ukey_DM(23 downto 16);
--         RAM(112) <= ukey_DM(31 downto 24);
     
          --Mode
--          RAM(136) <= x"00";
--          RAM(137) <= x"00";
--          RAM(138) <= x"00";
--          RAM(139) <= "0000" & mode_DM;
         
--          --Key Valid
--          RAM(144) <= x"00";
--          RAM(145) <= x"00";
--          RAM(146) <= x"00";
--          RAM(147) <= "0000000" & key_vld_DM;
      
       
       end if;
 end if;
 end process;
-- ram_addr <= mem_access_addr_DM(6 downto 0);
 
-- process(clk_DM, ram_addr, mem_write_en_DM, mem_write_data_DM)
--     begin
--      if(rising_edge(clk_DM)) then
--          if (mem_write_en_DM='1') then
--               ram(to_integer(unsigned(ram_addr)))   <= mem_write_data_DM(31 downto 24);
--               ram(to_integer(unsigned(ram_addr)+1)) <= mem_write_data_DM(23 downto 16);
--               ram(to_integer(unsigned(ram_addr)+2)) <= mem_write_data_DM(15 downto 8);
--               ram(to_integer(unsigned(ram_addr)+3)) <= mem_write_data_DM(7 downto 0);
--          end if;
--      end if;
-- end process;
   mem_read_data_DM <= ram(CONV_INTEGER(ram_addr)) & ram(CONV_INTEGER(ram_addr)+1) & 
                       ram(CONV_INTEGER(ram_addr)+2) & ram(CONV_INTEGER(ram_addr)+3) 
                       when (mem_read_DM='1') else x"00000000";


end Behavioral;