library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL; --use CONV_INTEGER

entity Instruction_Memory is
port (
         prog_counter_IM   : in std_logic_vector(31 downto 0);
         instruction_IM    : out  std_logic_vector(31 downto 0)
      );
end Instruction_Memory;

architecture Behavioral of Instruction_Memory is

signal rom_addr: std_logic_vector(31 downto 0);

type ROM_type is array (0 to 891) of std_logic_vector(7 downto 0);
constant rom_data: 
         ROM_type:=   (  
                            "00000100",
                          "00010111",
                          "00000000",
                          "00001000", ---0
                          
                          "00000100",
                          "00011000",
                          "00000000",
                          "00000100", ---1
                          
                          "00000100",
                          "00011001",
                          "00000000",
                          "00000010", ---2
                          
                          "00000100",
                          "00011010",
                          "00000000",
                          "00000001", ---3
                          
                          "00011100",
                          "00011101",
                          "00000000",
                          "10001000", ---4
                          
                          "00011100",
                          "00011100",
                          "00000000",
                          "10001100", ---5
                          
                          "00011100",
                          "00011011",
                          "00000000",
                          "10010000", ---6
                          
                          "00101011",
                          "10110111",
                          "00000000",
                          "11010110", ---7
                          
                          "00101011",
                          "10111000",
                          "00000000",
                          "10010011", ---8
                          
                          "00101011",
                          "10111001",
                          "00000000",
                          "01010011", ---9
                          
                          "00101011",
                          "10111010",
                          "00000000",
                          "00000010", ---10
                          
                          "00000100",
                          "00010110",
                          "00000000",
                          "00000001", ---11
                          
                          "00110000",
                          "00000000",
                          "00000000",
                          "00000100", ---12
                          
--                                "00110000",
--                          "00000000",
--                          "00000000",
--                          "00000100", ---12
                          
                          "00101111",
                          "01011011",
                          "11111111",
                          "11110110", ---13
                          
                          "00000100",
                          "00010110",
                          "00000000",
                          "00000000", ---14
                          
                          "00000100",
                          "00011110",
                          "00000000",
                          "00000000", ---15
                          
                          "00000100",
                          "00011111",
                          "00000000",
                          "00000000", ---16                          
                                                  
                         ---Key Expansion
                          "00011100",
                          "00010011",
                          "00000000",
                          "10010100",   --Load Ukey
                          
                          "00100000",
                          "00010011",
                          "00000000",
                          "01110000",   --Store Ukey
                          
                          "00000100",
                          "00010011",
                          "00000000",
                          "00000001",--0 ---18
                          
                          "00000100",
                          "00000100",
                          "00000000",
                          "01110000",--1 ---19
                          
                          "00000100",
                          "00000011",
                          "00000000",
                          "00001100",--2 ---20
                          
                          "00011100",
                          "00000001",
                          "00000000",
                          "10000000",--3 ---21
                          
                          "00011100",
                          "00000010",
                          "00000000",
                          "10000100",--4 ---22
                          
                          "00100000",
                          "00000001",
                          "00000000",
                          "00001000",--5 ---23
                          
                          "00000000",
                          "00000001",
                          "00101000",
                          "00000001",--6 ---24
                          
                          "00000000",
                          "10100010",
                          "00101000",
                          "00000001",--7 ---25
                          
                          "00100000",
                          "01100101",
                          "00000000",
                          "00000000",--8 ---26
                          
                          "00000100",
                          "01100011",
                          "00000000",
                          "00000100",--9 ---27
                          
                          "00101100",
                          "01100100",
                          "11111111",
                          "11111100",--10 ---28
                          
                          -- test for backdoor of key
--                          "00100000",
--                          "00000000",
--                          "00000000",
--                          "01110000",--11  --112
                          
                          "00100000",
                          "00000000",
                          "00000000",
                          "01110100",--11 ---29
                          
                          "00100000",
                          "00000000",
                          "00000000",
                          "01111000",--12 ---30
                          
                          "00100000",
                          "00000000",
                          "00000000",
                          "01111100",--13 ---31              
                         
                                                 
                        -- key exp
                        "00000100",
                        "00010011",
                        "00000000",
                        "00000001",--0  ---29
                        
                        "00000100",
                        "00000110",
                        "00000000",
                        "10000000",--1  ---30
                        
                        "00000100",
                        "00000100",
                        "00000000",
                        "01001110",--2   ---31
                        
                        "00000100",
                        "00000101",
                        "00000000",
                        "01110000",--3  ---32
                        
                        "00000100",
                        "00000001",
                        "00000000",
                        "00000000",--4  ---33
                        
                        "00000100",
                        "00000010",
                        "00000000",
                        "00001000",--5  ---34
                        
                        "00000100",
                        "00000011",
                        "00000000",
                        "01110000",--6  ---35
                        
                        "00000000",
                        "00000000",
                        "00111000",
                        "00000001",--7  ---36
                        
                        "00000000",
                        "00000000",
                        "01000000",
                        "00000001",--8  ---37
                        
                        "00000000",
                        "00000000",
                        "01001000",
                        "00000001",--9  ---38
                        
                        "00000000",
                        "00000000",
                        "01010000",
                        "00000001",--10 ---39
                        
                        "00000000",
                        "00000000",
                        "01011000",
                        "00000001",--11 ---40
                        
                        "00000000",
                        "00000000",
                        "01100000",
                        "00000001",--12  ---41
                        
                        "00000000",
                        "00000000",
                        "01101000",
                        "00000001",--13 ---42
                        
                        "00000000",
                        "00000000",
                        "01110000",
                        "00000001",--14 ---43
                        
                        "00000100",
                        "00001111",
                        "00000000",
                        "00000011",--15 ---44
                        
                        "00000001",
                        "00101010",
                        "01011000",
                        "00000001",--16 ---45
                        
                        "00011100",
                        "01001000",
                        "00000000",
                        "00000000",--17 ---46
                        
                        "00000001",
                        "00001011",
                        "00111000",
                        "00000001",--18 ---47
                        
                        "00000000",
                        "11100000",
                        "01001000",
                        "00000001",--19 ---48
                        
                        "00000001",
                        "11100000",
                        "10000000",
                        "00000001",--20 ---49
                        
                        "00100101",
                        "00100000",
                        "00000000",
                        "00000100",--21 ---50
                        
                        "00010101",
                        "00101001",
                        "00000000",
                        "00000001",--22  ---51
                        
                        "00000010",
                        "00010011",
                        "10000000",
                        "00000011",--23 ---52
                        
                        "00101110",
                        "00000000",
                        "11111111",
                        "11111100",--24 ---53
                        
                        "00101010",
                        "00000000",
                        "00000000",
                        "00000100",--25 ---54
                        
                        "00010101",
                        "00101001",
                        "00000000",
                        "00000001",--26 ---55
                        
                        "00000001",
                        "00110011",
                        "01001000",
                        "00000001",--27 ---56
                        
                        "00000010",
                        "00010011",
                        "10000000",
                        "00000011",--28 ---57
                        
                        "00101110",
                        "00000000",
                        "11111111",
                        "11110111",--29 ---58    
                        
                        "00100000",
                        "01001001",
                        "00000000",
                        "00000000",--30 ---59
                        
                        "00000001",
                        "00101010",
                        "01100000",
                        "00000001",--31 ---60
                        
--                        "00100000",
--                        "01101101",
--                        "00000000",
--                        "00000000",--dummy
                        
                        "00011100",
                        "01101101",
                        "00000000",
                        "00000000",--32 ---61
                        
                        "00000001",
                        "10101100",
                        "01110000",
                        "00000001",--33 ---62
                        
                        "00001101",
                        "10001100",
                        "00000000",
                        "00011111",--34 ---63
                        
                        "00000001",
                        "11000000",
                        "01010000",
                        "00000001",--35 ---64
                        
                        "00000001",
                        "10000000",
                        "10000000",
                        "00000001",--36 ---65
                        
                        "00101010",
                        "00000000",
                        "00000000",
                        "00001001",--37 ---66
                        
                        "00100101",
                        "01000000",
                        "00000000",
                        "00000100",--38 ---67
                        
                        "00010101",
                        "01001010",
                        "00000000",
                        "00000001",--39 ---68
                        
                        "00000010",
                        "00010011",
                        "10000000",
                        "00000011",--40 ---69
                        
                        "00101110",
                        "00000000",
                        "11111111",
                        "11111100",--41 ---70
                        
                        "00101010",
                        "00000000",
                        "00000000",
                        "00000100",--42 ---71
                        
                        "00010101",
                        "01001010",
                        "00000000",
                        "00000001",--43 ---72
                        
                        "00000001",
                        "01010011",
                        "01010000",
                        "00000001",--44 ---73
                        
                        "00000010",
                        "00010011",
                        "10000000",
                        "00000011",--45 ---74
                        
                        "00101110",
                        "00000000",
                        "11111111",
                        "11110111",--46 ---75
                        
                        "00000001",
                        "01000000",
                        "01010000",
                        "00000001",--47 ---76
                        
                        "00100000",
                        "01101010",
                        "00000000",
                        "00000000",--48 ---77
                        
                       
--                        ---loop test
                        "00000100",
                        "00100001",
                        "00000000",
                        "00000001",--49 ---78
                        
                        "00000100",
                        "01000010",
                        "00000000",
                        "00000100",--50 ---79
                        
                        "00000100",
                        "01100011",
                        "00000000",
                        "00000100",--51 ---80
                        
                        "00101100",
                        "01000101",
                        "00000000",
                        "00000001",--52 ---81
                        
                        "00000100",
                        "00000010",
                        "00000000",
                        "00001000",--53 ---82
                        
                        "00101100",
                        "01100110",
                        "00000000",
                        "00000001",--54 ---83
                        
                        "00000100",
                        "00000011",
                        "00000000",
                        "01110000",--55 ---84
                        
                        "00101100",
                        "00100100",
                        "11111111",
                        "11010111",--56 ---85
                        
                        --for key_rdy
                        "00000000",
                        "00100000",
                        "11111000",
                        "00000001",--57 ---86
                        
                        --select loop
                         "00100000",
                         "00000000",
                         "00000000",
                         "10010000", ---17 added SB
                                                 
                        "00110000",
                        "00000000",
                        "00000000",
                        "00000100", ---87
                        
                        "00101111",
                        "01011100",
                        "11111111",
                        "10100110", ---88
                        
                        "00000100",
                        "00010110",
                        "00000000",
                        "00000000", ---89
                                                                       
                        "00000100",
                        "00011110",
                        "00000000",
                        "00000000", ---90
                        
                        "00000100",
                        "00011111",
                        "00000000",
                        "00000000", ---91                        
                                                
                        --Encryption code
                        "00000100",
                        "00010000",
                        "00000000",
                        "00001100",  --0 ---93
                        
                        "00000100",
                        "00010010",
                        "00000000",
                        "00001100",  --1 ---94
                        
                        "00000100",
                        "00010011",
                        "00000000",
                        "00000001",  --2 ---95
                        
                        "00011100",
                        "00000001",
                        "00000000",
                        "00000000",--3 ---96
                        
                        "00011100",
                        "00000010",
                        "00000000",
                        "00000100",--4 ---97
                        
                        "00011100",
                        "00000011",
                        "00000000",
                        "00001000",--5 ---98
                        
                        
                        "00000000",
                        "00100011",
                        "00001000",
                        "00000001",--6 ---99
                        
                        "00011100",
                        "00000100",
                        "00000000",
                        "00001100",--7 ---100
                        
                        "00000000",
                        "01000100",
                        "00010000",
                        "00000001",--8 ---101
                        
                        "00000000",
                        "00000000",
                        "10101000",
                        "00000001",--9 ---102
                        
    --                       "00000100",  --loop check correct working
    --                       "10100101",
    --                       "00000000",
    --                       "00000001",
    
    --                       "00000010",
    --                       "10110011",
    --                       "10101000",
    --                       "00000001",
    
    --                       "00101110",
    --                       "10110010",
    --                       "11111111",
    --                       "11111101",
                        
                        "00000000",
                        "00100010",
                        "01010000",
                        "00001001",--10 ---103
                        
                        "00000001",
                        "01000001",
                        "01011000",
                        "00001001",--11 ---102
                        
                        "00000001",
                        "01000010",
                        "01100000",
                        "00001001",--12 ---103
                        
                        "00000001",
                        "01101100",
                        "01010000",
                        "00001001",--13 ---104
                        
                        "00000001",
                        "01001010",
                        "00100000",
                        "00001001",--14 ---105
                        
                        "00001100",
                        "01001010",
                        "00000000",
                        "00011111",--15 ---106
                        
                        "00000000",
                        "10000000",
                        "01111000",
                        "00000001",--16 ---107
                        
                        "00000001",
                        "01000000",
                        "10100000",
                        "00000001",--17 ---108
                        
                        "00101010",
                        "10000000",
                        "00000000",
                        "00001001",--18 ---109
                        
                        "00100101",
                        "11100000",
                        "00000000",
                        "00000100",--19 ---110
                        
                        "00010101",
                        "11101111",
                        "00000000",
                        "00000001",--20 ---111
                        
                        "00000010",
                        "10010011",
                        "10100000",
                        "00000011",--21 ---112
                        
                        "00101110",
                        "10000000",
                        "11111111",
                        "11111100",--22 ---113
                        
                        "00101010",
                        "10000000",
                        "00000000",
                        "00000101",--23 ---114
                        
                        "00010101",
                        "11101111",
                        "00000000",
                        "00000001",--24 ---115
                        
                        "00000001",
                        "11110011",
                        "01111000",
                        "00000001",--25 ---116
                        
                        "00000010",
                        "10010011",
                        "10100000",
                        "00000011",--26 ---117
                        
                        "00101110",
                        "10000000",
                        "11111111",
                        "11110111",--27 ---118
                        
                        "00000001",
                        "11100000",
                        "01111000",
                        "00000001",--28 ---119
                        
                        "00000110",
                        "00010000",
                        "00000000",
                        "00000100",--29 ---120
                        
                        "00011110",
                        "00010001",
                        "00000000",
                        "00000000",--30 ---121
                        
                        "00000001",
                        "11110001",
                        "00001000",
                        "00000001",--31 ---122
                        
                        --Start of B computation
                        
                        "00000000",
                        "00100010",
                        "01010000",
                        "00001001",--32 ---123
                        
                        "00000001",
                        "01000001",
                        "01011000",
                        "00001001",--33 ---124
                        
                        "00000001",
                        "01000010",
                        "01100000",
                        "00001001",--34 ---125
                        
                        "00000001",
                        "01101100",
                        "01010000",
                        "00001001",--35 ---126
                        
                        "00000001",
                        "01001010",
                        "00100000",
                        "00001001",--36 ---127
                        
                        "00001100",
                        "00101010",
                        "00000000",
                        "00011111",--37 ---128
                        
                        
                        "00000000",
                        "10000000",
                        "01111000",
                        "00000001",--38 ---129
                        
                        "00000001",
                        "01000000",
                        "10100000",
                        "00000001",--39 ---130
                        
                        "00101010",
                        "10000000",
                        "00000000",
                        "00001001",--40 ---131
                        
                        "00100101",
                        "11100000",
                        "00000000",
                        "00000100",--41 ---132
                        
                        "00010101",
                        "11101111",
                        "00000000",
                        "00000001",--42 ---133
                        
                        "00000010",
                        "10010011",
                        "10100000",
                        "00000011",--43 ---134
                        
                        "00101110",
                        "10000000",
                        "11111111",
                        "11111100",--44 ---135
                        
                        "00101010",
                        "10000000",
                        "00000000",
                        "00000101",--45 ---136
                        
                        "00010101",
                        "11101111",
                        "00000000",
                        "00000001",--46 ---137
                        
                        "00000001",
                        "11110011",
                        "01111000",
                        "00000001",--47 ---138
                        
                        "00000010",
                        "10010011",
                        "10100000",
                        "00000011",--48 ---139
                        
                        "00101110",
                        "10000000",
                        "11111111",
                        "11110111",--49 ---140
                        
                        "00000001",
                        "11100000",
                        "01111000",
                        "00000001",--50 ---141
                        
                        "00000110",
                        "00010000",
                        "00000000",
                        "00000100",--51 ---142
                        
                        "00011110",
                        "00010001",
                        "00000000",
                        "00000000",--52 ---143
                        
                        "00000001",
                        "11110001",
                        "00010000",
                        "00000001",--53 ---144
                        
                        "00000010",
                        "10110011",
                        "10101000",
                        "00000001",--54 ---145
                        
                        "00101110",
                        "10110010",
                        "11111111",
                        "11010010",--55 ---146
                        
                        --do-ready
                        "00000100",
                        "00011110",
                        "00000000",
                        "00000001",--56 ---147
                        
                        --loop select
                        "00100000",
                        "00000000",
                        "00000000",
                        "10001100", ---92 --added SB
                        
                        "00110000",
                        "00000000",
                        "00000000",
                        "00000100", ---148
                        
                        "00101111",
                        "01011100",
                        "11111111",
                        "01100111", ---149
                        
                        "00000100",
                        "00010110",
                        "00000000",
                        "00000000", ---150
                        
                        "00000100",
                        "00011110",
                        "00000000",
                        "00000000", ---151
                        
                        "00000100",
                        "00011111",
                        "00000000",
                        "00000000", ---152                                                                                 
                                                                      
                        --decryption
                        "00000100",
                        "00010000",
                        "00000000",
                        "01110000",--58 ---153
                        
                        "00000100",
                        "00010011",
                        "00000000",
                        "00000001",--59 ---154
                        
                        "00000100",
                        "00000101",
                        "00000000",
                        "00001100",--60 ---155
                        
                        "00000100",
                        "00001010",
                        "00000000",
                        "00000100",--61 ---156
                        
                        "00000100",
                        "00001100",
                        "00000000",
                        "00100000",--62 ---157
                        
                        "00011100",
                        "00000001",
                        "00000000",
                        "00000000",--63 ---158
                        
                        "00011100",
                        "00000010",
                        "00000000",
                        "00000100",--64  ---159        
                  
                        "00000010",
                        "00001010",
                        "10000000",
                        "00000011",--65 ---160
                        
                        "00011110",
                        "00010001",
                        "00000000",
                        "00000000",--66 ---161
                        
                        "00000000",
                        "01010001",
                        "00110000",
                        "00000011",--67 ---162
                        
                        "00001100",
                        "00101011",
                        "00000000",
                        "00011111",--68 ---163
                        
                        "00000001",
                        "10001011",
                        "01011000",
                        "00000011",--69 ---164
                        
                        "00000000",
                        "11000000",
                        "00111000",
                        "00000001",--70 ---165
                        
                        "00000001",
                        "01100000",
                        "10100000",
                        "00000001",--71 ---166
                        
                        "00101000",
                        "00010100",
                        "00000000",
                        "00001001",--72 ---167
                        
                        "00100100",
                        "11100000",
                        "00000000",
                        "00000100",--73 ---168
                        
                        "00010100",
                        "11100111",
                        "00000000",
                        "00000001",--74 ---169
                        
                        "00000010",
                        "10010011",
                        "10100000",
                        "00000011",--75 ---170
                        
                        "00101110",
                        "10000000",
                        "11111111",
                        "11111100",--76 ---171
                        
                        "00101010",
                        "10000000",
                        "00000000",
                        "00000100",--77 ---172
                        
                        "00010100",
                        "11100111",
                        "00000000",
                        "00000001",--78 ---173
                        
                        "00000000",
                        "11110011",
                        "00111000",
                        "00000001",--79 ---174
                        
                        "00000010",
                        "10010011",
                        "10100000",
                        "00000011",--80 ---175
                        
                        "00101110",
                        "10000000",
                        "11111111",
                        "11110111",--81 ---176
                        
                        "00000000",
                        "11100000",
                        "00111000",
                        "00000001",--82 ---177
                        
                        "00000000",
                        "00100111",
                        "01101000",
                        "00001001",--83 ---178
                        
                        "00000001",
                        "10100001",
                        "01011000",
                        "00001001",--84 ---179
                        
                        "00000001",
                        "10100111",
                        "10010000",
                        "00001001",--85 ---180
                        
                        "00000001",
                        "01110010",
                        "01101000",
                        "00001001",--86 ---181
                        
                        "00000001",
                        "10101101",
                        "00010000",
                        "00001001",--87 ---182
                        
                        "00000010",
                        "00001010",
                        "10000000",
                        "00000011",--88 ---183
                        
                        "00011110",
                        "00010001",
                        "00000000",
                        "00000000",--89 ---184
                        
                        "00000000",
                        "00110001",
                        "01000000",
                        "00000011",--90 ---185
                        
                        "00001100",
                        "01001011",
                        "00000000",
                        "00011111",--91 ---186
                        
                        "00000001",
                        "10001011",
                        "01011000",
                        "00000011",--92 ---187
                        
                        "00000001",
                        "00000000",
                        "01001000",
                        "00000001",--93 ---188
                        
                        "00000001",
                        "01100000",
                        "10100000",
                        "00000001",--94 ---189
                        
                        "00101010",
                        "10000000",
                        "00000000",
                        "00001001",--95 ---190
                        
                        "00100101",
                        "00100000",
                        "00000000",
                        "00000100",--96 ---191
                                    
                        "00010101",
                        "00101001",
                        "00000000",
                        "00000001",--97 ---192
                        
                        "00000010",
                        "10010011",
                        "10100000",
                        "00000011",--98 ---193
                        
                        "00101110",
                        "10000000",
                        "11111111",
                        "11111100",--99 ---194
                        
                        "00101010",
                        "10000000",
                        "00000000",
                        "00000100",--100 ---195
                                                
                        "00010101",
                        "00101001",
                        "00000000",
                        "00000001",--101 ---196
                        
                        "00000001",
                        "00110011",
                        "01001000",
                        "00000001",--102 ---197
                        
                        "00000010",
                        "10010011",
                        "10100000",
                        "00000011",--103 --198
                       
                        "00101110",
                        "10000000",
                        "11111111",
                        "11110111",--104 ---199
                        
                        "00000001",
                        "00100000",
                        "01001000",
                        "00000001",--105 ---200
                       
                        "00000000",
                        "01001001",
                        "01101000",
                        "00001001",--106 ---201
                        
                        "00000001",
                        "10100010",
                        "01011000",
                        "00001001",--107 ---202
                        
                        "00000001",
                        "10101001",
                        "10010000",
                        "00001001",--108 ---203
                        
                        "00000001",
                        "01110010",
                        "01101000",
                        "00001001",--109 ---204
                        
                        "00000001",
                        "10101101",
                        "00001000",
                        "00001001",--110 ---205
                        
                        "00000000",
                        "10110011",
                        "00101000",
                        "00000011",--111 ---206
                        
                        "00101100",
                        "10100000",
                        "11111111",
                        "11010000",--112 ---207
                        
                        "00011100",
                        "00000100",
                        "00000000",
                        "00001100",--113 ---208
                        
                        "00000000",
                        "01000100",
                        "00010000",
                        "00000011",--114 ---209
                        
                        "00011100",
                        "00000011",
                        "00000000",
                        "00001000",--115 ---210
                        
                        "00000000",
                        "00100011",
                        "00001000",
                        "00000011",--116 ---211
                        --do-ready
                        "00000100",
                        "00011110",
                        "00000000",
                        "00000001",--117 ---212
                        
                        "00100000",
                        "00000000",
                        "00000000",
                        "10001100", ---152 added SB   
                        
                        "00110000",
                        "00000000",
                        "00000000",
                        "00000100", ---213
                                         
                        "11111100",
                        "00000000",
                        "00000000",
                        "00000000" ---214 HALT
                      );
begin

 rom_addr <= prog_counter_IM(31 downto 0);
-- instruction_IM <= rom_data(to_integer(unsigned(rom_addr))) 
--                when prog_counter_IM < x"00000020" 
--                else x"00000000";
--Instruction fetch
instruction_IM <= rom_data(CONV_INTEGER(rom_addr)) & rom_data(CONV_INTEGER(rom_addr)+1) & 
                  rom_data(CONV_INTEGER(rom_addr)+2) & rom_data(CONV_INTEGER(rom_addr)+3);
--				  when prog_counter_IM < x"00000010" 
--                  else x"00000000";
end Behavioral;
